//Byte level FSM commands
`define START 'b100
`define STOP 'b101
`define RWACK 'b010
`define RWNACK 'b011
`define WRITE 'b001
`define SETBUS 'b110
`define WAIT 'b000

//Register blocks
`define CSR 'b00
`define DPR 'b01
`define CMDR 'b10
`define FSMR 'b11

